module ALU(
    input logic [1:0] a, b,
    input logic select,
    output logic [1:0] out
):


endmodule